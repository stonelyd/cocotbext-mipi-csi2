/*
 * Basic CSI-2 test module
 *
 * Copyright (c) 2024 CSI-2 Extension Contributors
 */

`timescale 1ns / 1ps

module test_csi2_basic (
    input  wire clk,
    input  wire reset_n,

    // D-PHY Clock Lane
    output wire clk_p,
    output wire clk_n,

    // D-PHY Data Lane 0
    output wire data0_p,
    output wire data0_n,

    // D-PHY Data Lane 1 (for multi-lane tests)
    output wire data1_p,
    output wire data1_n,

    // Status signals
    output reg  frame_valid,
    output reg  line_valid,
    output reg [7:0] pixel_data,
    output reg  pixel_valid
);

    // Simple CSI-2 receiver implementation for testing
    // This is a minimal implementation to validate the TX model

    reg [3:0] state;
    reg [7:0] byte_buffer;
    reg [2:0] bit_count;
    reg [15:0] packet_length;
    reg [15:0] byte_count;

    // State machine states
    localparam IDLE = 4'h0;
    localparam HS_SYNC = 4'h1;
    localparam HEADER = 4'h2;
    localparam PAYLOAD = 4'h3;
    localparam CHECKSUM = 4'h4;

    // Decode differential signals (simplified)
    wire clk_lane = clk_p & ~clk_n;
    wire data0_lane = data0_p & ~data0_n;
    wire data1_lane = data1_p & ~data1_n;

    // Packet header fields
    reg [7:0] data_id;
    reg [15:0] word_count;
    reg [7:0] ecc;

    // Virtual channel and data type
    wire [1:0] virtual_channel = data_id[7:6];
    wire [5:0] data_type = data_id[5:0];

    // Frame and line tracking
    reg frame_active;
    reg line_active;
    reg [15:0] current_frame;
    reg [15:0] current_line;

    always @(posedge clk) begin
        if (!reset_n) begin
            state <= IDLE;
            frame_valid <= 1'b0;
            line_valid <= 1'b0;
            pixel_valid <= 1'b0;
            pixel_data <= 8'h00;
            byte_buffer <= 8'h00;
            bit_count <= 3'h0;
            packet_length <= 16'h0;
            byte_count <= 16'h0;
            frame_active <= 1'b0;
            line_active <= 1'b0;
            current_frame <= 16'h0;
            current_line <= 16'h0;
        end else begin
            case (state)
                IDLE: begin
                    // Wait for HS sync pattern
                    if (data0_lane) begin
                        state <= HS_SYNC;
                        bit_count <= 3'h0;
                    end
                end

                HS_SYNC: begin
                    // Accumulate bits into bytes
                    byte_buffer <= {data0_lane, byte_buffer[7:1]};
                    bit_count <= bit_count + 1;

                    if (bit_count == 7) begin
                        // Complete byte received
                        if (byte_count < 4) begin
                            // Header bytes
                            case (byte_count)
                                0: data_id <= {data0_lane, byte_buffer[7:1]};
                                1: word_count[7:0] <= {data0_lane, byte_buffer[7:1]};
                                2: word_count[15:8] <= {data0_lane, byte_buffer[7:1]};
                                3: ecc <= {data0_lane, byte_buffer[7:1]};
                            endcase
                            byte_count <= byte_count + 1;

                            if (byte_count == 3) begin
                                // Header complete
                                packet_length <= word_count;
                                if (word_count == 0) begin
                                    // Short packet
                                    state <= IDLE;
                                    process_short_packet();
                                end else begin
                                    // Long packet
                                    state <= PAYLOAD;
                                end
                                byte_count <= 0;
                            end
                        end
                        bit_count <= 0;
                        byte_buffer <= 0;
                    end
                end

                PAYLOAD: begin
                    // Receive payload data
                    byte_buffer <= {data0_lane, byte_buffer[7:1]};
                    bit_count <= bit_count + 1;

                    if (bit_count == 7) begin
                        // Complete payload byte
                        pixel_data <= {data0_lane, byte_buffer[7:1]};
                        pixel_valid <= 1'b1;

                        byte_count <= byte_count + 1;
                        if (byte_count >= packet_length - 1) begin
                            state <= CHECKSUM;
                            byte_count <= 0;
                        end

                        bit_count <= 0;
                        byte_buffer <= 0;
                    end else begin
                        pixel_valid <= 1'b0;
                    end
                end

                CHECKSUM: begin
                    // Receive checksum (2 bytes)
                    byte_buffer <= {data0_lane, byte_buffer[7:1]};
                    bit_count <= bit_count + 1;

                    if (bit_count == 7) begin
                        byte_count <= byte_count + 1;
                        if (byte_count >= 1) begin
                            // Packet complete
                            state <= IDLE;
                            byte_count <= 0;
                        end
                        bit_count <= 0;
                        byte_buffer <= 0;
                    end
                end
            endcase
        end
    end

    // Process short packets
    task process_short_packet;
        begin
            case (data_type)
                6'h00: begin // Frame Start
                    frame_active <= 1'b1;
                    frame_valid <= 1'b1;
                    current_frame <= word_count;
                    $display("Frame Start: VC=%d, Frame=%d", virtual_channel, word_count);
                end

                6'h01: begin // Frame End
                    frame_active <= 1'b0;
                    frame_valid <= 1'b0;
                    line_active <= 1'b0;
                    line_valid <= 1'b0;
                    $display("Frame End: VC=%d, Frame=%d", virtual_channel, word_count);
                end

                6'h02: begin // Line Start
                    line_active <= 1'b1;
                    line_valid <= 1'b1;
                    current_line <= word_count;
                    $display("Line Start: VC=%d, Line=%d", virtual_channel, word_count);
                end

                6'h03: begin // Line End
                    line_active <= 1'b0;
                    line_valid <= 1'b0;
                    $display("Line End: VC=%d, Line=%d", virtual_channel, word_count);
                end

                6'h08, 6'h09, 6'h0A, 6'h0B, 6'h0C, 6'h0D, 6'h0E, 6'h0F: begin // Generic Short Packets
                    $display("Generic Short Packet: DT=0x%02x, VC=%d, Data=0x%04x",
                            data_type, virtual_channel, word_count);
                end

                6'h18, 6'h19, 6'h1A, 6'h1C, 6'h1D, 6'h1E, 6'h1F: begin // YUV Data Types
                    $display("YUV Data Packet: DT=0x%02x, VC=%d, Data=0x%04x",
                            data_type, virtual_channel, word_count);
                end

                6'h20, 6'h21, 6'h22, 6'h23, 6'h24: begin // RGB Data Types
                    $display("RGB Data Packet: DT=0x%02x, VC=%d, Data=0x%04x",
                            data_type, virtual_channel, word_count);
                end

                6'h28, 6'h29, 6'h2A, 6'h2B, 6'h2C, 6'h2D, 6'h2E, 6'h2F: begin // RAW Data Types
                    $display("RAW Data Packet: DT=0x%02x, VC=%d, Data=0x%04x",
                            data_type, virtual_channel, word_count);
                end

                6'h30, 6'h31, 6'h32, 6'h33, 6'h34, 6'h35, 6'h36, 6'h37: begin // User Defined Types
                    $display("User Defined Packet: DT=0x%02x, VC=%d, Data=0x%04x",
                            data_type, virtual_channel, word_count);
                end

                default: begin
                    $display("Unknown short packet: DT=0x%02x, VC=%d, Data=0x%04x",
                            data_type, virtual_channel, word_count);
                end
            endcase
        end
    endtask

    // Generate differential clock (simplified)
    reg clk_out;
    always @(posedge clk) begin
        if (reset_n) begin
            clk_out <= ~clk_out;
        end else begin
            clk_out <= 1'b0;
        end
    end

    assign clk_p = clk_out;
    assign clk_n = ~clk_out;

    // Initially tri-state data lanes
    assign data0_p = 1'bz;
    assign data0_n = 1'bz;
    assign data1_p = 1'bz;
    assign data1_n = 1'bz;

endmodule
